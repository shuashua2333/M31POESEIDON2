`timescale 1ns/1ps
package m31_constants_pkg;
    import m31_pkg::*;

    // Define a packed state type for WIDTH=16
    typedef m31_t [15:0] state16_t;

    // Initial Round Constants (Added before S-box)
    // Format: ROUND_CONSTS_INITIAL[round_idx] returns a packed array of 16 elements
    localparam state16_t ROUND_CONSTS_INITIAL [0:3] = '{
        '{31'd1614794869, 31'd733565087, 31'd1248974626, 31'd1395707998, 31'd1606546523, 31'd308743513, 31'd933669702, 31'd1509218160, 31'd857651441, 31'd974826695, 31'd1777538858, 31'd1732216065, 31'd1121120522, 31'd867595173, 31'd2052960689, 31'd670752198},
        '{31'd354722588, 31'd553962986, 31'd836569592, 31'd974777474, 31'd478426997, 31'd1010294888, 31'd1451694789, 31'd1745808542, 31'd1022914986, 31'd615368408, 31'd358422393, 31'd1563765150, 31'd1735187654, 31'd2055660101, 31'd311580733, 31'd1457687568},
        '{31'd107763776, 31'd968153742, 31'd1642480066, 31'd1781773041, 31'd1610545562, 31'd2100202195, 31'd365270850, 31'd821769216, 31'd743793854, 31'd1777322674, 31'd511348931, 31'd1575313895, 31'd1314307614, 31'd1171073730, 31'd957403621, 31'd1099724285},
        '{31'd1609172128, 31'd1281424936, 31'd1121275927, 31'd1538050768, 31'd934311777, 31'd1656304581, 31'd1491107118, 31'd695522824, 31'd1017368981, 31'd1347088819, 31'd372969254, 31'd699322108, 31'd1825005418, 31'd670079580, 31'd1048805912, 31'd304102504}
    };

    // Internal Round Constants (Added to first element only)
    localparam m31_t ROUND_CONSTS_INTERNAL [0:13] = '{
        31'd129024239, 31'd1282387121, 31'd2004475442, 31'd535738304, 31'd1985680653, 31'd895998816, 31'd1108547306, 31'd776893336, 31'd1108245527, 31'd574331301, 31'd1825109420, 31'd1194870642, 31'd1497066195, 31'd1664793266
    };

    // Terminal Round Constants
    localparam state16_t ROUND_CONSTS_TERMINAL [0:3] = '{
        '{31'd2135403312, 31'd1833171446, 31'd1217130568, 31'd1610027373, 31'd437172020, 31'd2020259742, 31'd2143547951, 31'd802809388, 31'd122792040, 31'd151742200, 31'd1491417545, 31'd359041126, 31'd802016690, 31'd16103019, 31'd2055094098, 31'd302658704},
        '{31'd848039704, 31'd1735444335, 31'd1574838747, 31'd1536582683, 31'd1943893587, 31'd718747682, 31'd4549961, 31'd367271168, 31'd696367131, 31'd1495214374, 31'd458819359, 31'd1766051075, 31'd2058149815, 31'd1580136315, 31'd173288461, 31'd60728125},
        '{31'd1183379851, 31'd1790329919, 31'd2117379525, 31'd37211066, 31'd1687696498, 31'd618979668, 31'd1160504957, 31'd297763826, 31'd1082619536, 31'd1744615017, 31'd782638163, 31'd2077368442, 31'd1004172913, 31'd427470023, 31'd173154748, 31'd1689611743},
        '{31'd688337540, 31'd1667233644, 31'd210718841, 31'd926128391, 31'd1823128363, 31'd1722126248, 31'd1214340530, 31'd637696247, 31'd95801870, 31'd1929310598, 31'd1903150401, 31'd1080767281, 31'd1927785244, 31'd723170958, 31'd1229207547, 31'd545339302}
    };
endpackage
